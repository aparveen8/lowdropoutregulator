* c:\users\aparv\esim-workspace\ayesha_LDO\ayesha_LDO.cir 
.lib "C:\FOSSEE\eSim\library\sky130_fd_pr\models\sky130.lib.spice" tt 

******* Transistor Connection*****
xMN4   net_d    vbias2     net3     GND  sky130_fd_pr__nfet_01v8
xMP2   net1     net_d   VDD      VDD  sky130_fd_pr__pfet_01v8
xMN1   net3     VFB  net_diff GND  sky130_fd_pr__nfet_01v8
xM4  Vpass   vbias2     net4     GND  sky130_fd_pr__nfet_01v8
xM1  net4     VREF    net_diff GND  sky130_fd_pr__nfet_01v8
xMP3   net_d    vbias1     net1     VDD  sky130_fd_pr__pfet_01v8
xM3  Vpass   vbias1     net2     VDD  sky130_fd_pr__pfet_01v8
xMn5  net_diff VDD     GND      GND  sky130_fd_pr__nfet_01v8
xM5   VDD      VDD     GND      GND  sky130_fd_pr__nfet_01v8
xMP1  Vreg     Vpass  VDD      VDD  sky130_fd_pr__pfet_01v8
xMV2  net2     net_d   VDD      VDD  sky130_fd_pr__pfet_01v8
CL    Vreg     GND     10p
cc Vpass Vreg 1p

* Feedback resistors
RFB1   Vreg     VFB    150k
RFB2   VFB   GND       600k

***** Power *******

* Define Vdd as PWL for line transient response
Vdd vdd 0 PWL(0 1.5 1n 1.5 1.01n 2.5 2n 2.5 2.01n 1.8 3n 1.8 3.01n 3)
Vbias1 vbias1 0 0
vbias2 vbias2 0 3.3
VREF VREF 0 1.2

**** Analysis*****

* Perform transient analysis over a range that covers the PWL steps
.tran 0.1n 5n

* Control Statements

.control
run

**** Output Plot****

* Plot Vreg to observe the LDO's regulation response to Vdd variations
plot V(vdd) V(Vreg)

.endc
.end
